/*-----------------------------------------------------------------
File name     : yapp_tx_seqs.sv
Developers    : Kathleen Meade, Brian Dickinson
Created       : 01/04/11
Description   : YAPP UVC simple TX test sequence for labs 2 to 4
Notes         : From the Cadence "SystemVerilog Advanced Verification with UVM" training
-------------------------------------------------------------------
Copyright Cadence Design Systems (c)2015
-----------------------------------------------------------------*/

//------------------------------------------------------------------------------
//
// SEQUENCE: base yapp sequence - base sequence with objections from which 
// all sequences can be derived
//
//------------------------------------------------------------------------------
class yapp_base_seq extends uvm_sequence #(yapp_packet);
  
  // Required macro for sequences automation
  `uvm_object_utils(yapp_base_seq)

  // Constructor
  function new(string name="yapp_base_seq");
    super.new(name);
  endfunction

  task pre_body();
    uvm_phase phase;
    `ifdef UVM_VERSION_1_2
      // in UVM1.2, get starting phase from method
      phase = get_starting_phase();
    `else
      phase = starting_phase;
    `endif
    if (phase != null) begin
      phase.raise_objection(this, get_type_name());
      `uvm_info(get_type_name(), "raise objection", UVM_MEDIUM)
    end
  endtask : pre_body

  task post_body();
    uvm_phase phase;
    `ifdef UVM_VERSION_1_2
      // in UVM1.2, get starting phase from method
      phase = get_starting_phase();
    `else
      phase = starting_phase;
    `endif
    if (phase != null) begin
      phase.drop_objection(this, get_type_name());
      `uvm_info(get_type_name(), "drop objection", UVM_MEDIUM)
    end
  endtask : post_body

endclass : yapp_base_seq

//------------------------------------------------------------------------------
//
// SEQUENCE: yapp_5_packets
//
//  Configuration setting for this sequence
//    - update <path> to be hierarchial path to sequencer 
//
//  uvm_config_wrapper::set(this, "<path>.run_phase",
//                                 "default_sequence",
//                                 yapp_5_packets::get_type());
//
//------------------------------------------------------------------------------
class yapp_5_packets extends yapp_base_seq;
  
  // Required macro for sequences automation
  `uvm_object_utils(yapp_5_packets)

  // Constructor
  function new(string name="yapp_5_packets");
    super.new(name);
  endfunction

  // Sequence body definition
  virtual task body();
    `uvm_info(get_type_name(), "Executing yapp_5_packets sequence", UVM_LOW)
     repeat(5)
      `uvm_do(req)
  endtask
  
endclass : yapp_5_packets


class yapp_1_seq extends yapp_base_seq;

  `uvm_object_utils(yapp_1_seq)

  function new(string name="yapp_1_seq");
    super.new(name);
  endfunction

  task body();
    `uvm_info("SEQ", "yapp_1_seq", UVM_LOW)
    `uvm_do_with(req, {req.addr == 1;})
  endtask

endclass : yapp_1_seq


class yapp_012_seq extends yapp_base_seq;

  `uvm_object_utils(yapp_012_seq)

  function new(string name="yapp_012_seq");
    super.new(name);
  endfunction

  task body();
    `uvm_info("SEQ", "yapp_012_seq", UVM_LOW)
    `uvm_do_with(req, {req.addr == 0;})
    `uvm_do_with(req, {req.addr == 1;})
    `uvm_do_with(req, {req.addr == 2;})
  endtask

endclass : yapp_012_seq


class yapp_111_seq extends yapp_base_seq;

  `uvm_object_utils(yapp_111_seq)

  yapp_1_seq y1s;

  function new(string name="yapp_111_seq");
    super.new(name);
  endfunction

  task body();
    `uvm_info("SEQ", "yapp_111_seq", UVM_LOW)
    `uvm_do(y1s)
    `uvm_do(y1s)
    `uvm_do(y1s)
  endtask

endclass : yapp_111_seq


class yapp_repeat_addr_seq extends yapp_base_seq;

  `uvm_object_utils(yapp_repeat_addr_seq)

  rand logic [1:0] repeat_addr;

  constraint addr_c {repeat_addr != 3;}

  function new(string name="yapp_repeat_addr_seq");
    super.new(name);
  endfunction

  task body();
    `uvm_info("SEQ", "yapp_repeat_addr_seq", UVM_LOW)
    `uvm_do_with(req, {req.addr == repeat_addr;})
    `uvm_do_with(req, {req.addr == repeat_addr;})
  endtask

endclass : yapp_repeat_addr_seq


class yapp_incr_payload_seq extends yapp_base_seq;

  `uvm_object_utils(yapp_incr_payload_seq)

  function new(string name="yapp_incr_payload_seq");
    super.new(name);
  endfunction

  task body();
    `uvm_info("SEQ", "yapp_incr_payload_seq", UVM_LOW)
    `uvm_create(req)
    if (!req.randomize()) begin
    `uvm_error("RAND_FAIL", "Randomization of y1s packet failed")
    end
    foreach(req.payload[i]) begin
      req.payload[i] = i;
    end
    req.set_parity();
    `uvm_send(req)
  endtask

endclass : yapp_incr_payload_seq


class yapp_exhaustive_seq extends yapp_base_seq;

  `uvm_object_utils(yapp_exhaustive_seq)

  yapp_1_seq y1s;
  yapp_012_seq y012s;
  yapp_111_seq y111s;
  yapp_repeat_addr_seq yreps;
  yapp_incr_payload_seq yincs;

  function new(string name="yapp_exhaustive_seq");
    super.new(name);
  endfunction

  task body();
    `uvm_info("SEQ", "yapp_exhaustive_seq", UVM_LOW)
    `uvm_do(y1s)
    `uvm_do(y012s)
    `uvm_do(y111s)
    `uvm_do(yreps)
    `uvm_do(yincs)
  endtask

endclass : yapp_exhaustive_seq